module imem(input logic[5:0] a,
            output logic[31:0]rd);


logic[31:0] RAM[0:20] = {
    // ========== 阶段1：初始化（无冲突，确保值正确） ==========
    32'h2002000A,  // RAM[0]：addi $2, $0, 10  → $2=10（out[0]）
    32'h20030003,  // RAM[1]：addi $3, $0, 3   → $3=3（out[1]）
    32'h20040000,  // RAM[2]：addi $4, $0, 0   → $4=0（out[2]）
    32'h20050000,  // RAM[3]：addi $5, $0, 0   → $5=0（out[3]）
    32'h20070050,  // RAM[4]：addi $7, $0, 80  → $7=80（jr跳转至RAM[20]，80/4=20）
    
    // ========== 阶段2：基础R型指令 ==========
    32'h00431020,  // RAM[5]：add $2, $2, $3   → $2=10+3=13
    32'h00431822,  // RAM[6]：sub $3, $2, $3   → $3=13-3=10
    32'h00432024,  // RAM[7]：and $4, $2, $3   → $4=13&10=8
    32'h00432825,  // RAM[8]：or  $5, $2, $3   → $5=13|10=15
    32'h00852026,  // RAM[9]：xor $4, $4, $5   → $4=8^15=7
    32'h0043382A,  // RAM[10]：slt $7, $2, $3  → $7=0（13<10不成立）
    
    // ========== 阶段3：I型逻辑指令 ==========
    32'h3044000F,  // RAM[11]：andi $4, $2, 15 → $4=13&15=13
    32'h3465000F,  // RAM[12]：ori $5, $3, 15  → $5=10|15=15
    
    // ========== 阶段4：访存指令（简化，无冲突） ==========
    32'hAC020000,  // RAM[13]：sw $2, 0($0)    → 存储$2=13到地址0
    32'h8C030000,  // RAM[14]：lw $3, 0($0)    → 加载13到$3
    
    // ========== 阶段5：分支指令（修正偏移量） ==========
    32'h10430001,  // RAM[15]：beq $2,$3,1     → 偏移量1，跳转至RAM[17]（正确计算）
    32'h14470000,  // RAM[16]：bne $2,$7,0     → $2=13≠$7=0，不跳转
    32'h20420001,  // RAM[17]：addi $2, $2, 1  → $2=14（跳转后执行）
    
    // ========== 阶段6：jr跳转（修正地址，多跳3行） ==========
    32'h20070050,  // RAM[18]：addi $7, $0, 80 → $7=80（RAM[20]=80/4=20）
    32'h00E00008,  // RAM[19]：jr $7          → 跳转到RAM[20]（多跳1行，无越界）
    32'h00000000   // RAM[20]：nop            → 程序正常结束
};

// 超出指令范围返回空指令（nop），避免不定态
// 注意：流水线设计会使得程序最后重复返回自身(0x1000ffff)不可行
assign rd = (a <= 20) ? RAM[a] : 32'h00000000;
endmodule